module dec2bin( output )